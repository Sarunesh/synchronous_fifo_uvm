class sync_fifo_rd_seq extends uvm_sequence#(sync_fifo_rd_seq_item);
	//Factory registration
	`uvm_object_utils(sync_fifo_rd_seq)

	//Constructor
	`NEW_OBJECT
endclass: sync_fifo_rd_seq
