typedef uvm_sequencer#(sync_fifo_wr_seq_item) sync_fifo_wr_sqr;
