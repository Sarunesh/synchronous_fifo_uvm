class sync_fifo_rd_sqr extends uvm_sequencer#(sync_fifo_rd_seq_item);
//Factory registration
	`uvm_component_utils(sync_fifo_rd_sqr)
//Constructor
	`NEW_COMPONENT
endclass: sync_fifo_rd_sqr
