class sync_fifo_wr_sqr extends uvm_sequencer#(sync_fifo_wr_seq_item);
//Factory registration
	`uvm_component_utils(sync_fifo_wr_sqr)
//Constructor
	`NEW_COMPONENT
endclass: sync_fifo_wr_sqr
