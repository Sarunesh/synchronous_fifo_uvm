typedef uvm_sequencer#(sync_fifo_rd_seq_item) sync_fifo_rd_sqr;
